`include "pipeline.svh"
module mmu(
    
);
    
endmodule